
/* or.v */


module or_m (
    input       a, b,
    output wire c
);

    assign c = a | b;

endmodule
